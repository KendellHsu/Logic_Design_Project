module draw_main_scene (
    input clk,
    input rst,
    input [1:0] current_state, // Current game state
    input [1:0] selected_song,  // Selected song
    output reg [6143:0] menuMap  // Output to RGB matrix
);

    // State encoding
    localparam START_SCENE = 2'b00;
    localparam SONG_SELECT = 2'b01;
    localparam GAME_PLAY = 2'b10;
    localparam GAME_OVER = 2'b11;

    // Toggle for animation
    reg toggle;
    reg [20:0] counter;
    localparam animation_fps = 20'd160000;

    // Map definitions for different screens
    localparam start_scene_map_off = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111101101110110110110110110101101101110110101101101110110110110110110101101110110110110101101110110101101110110101101110110110110110101110110110110110110101110101101101110110101101101111000000111101101110110110110110110000101110000000110101101110110110110110110000110110000000110110101110110000101110110000101110110110110000000110110110110110110000110110101101110110000101101111000000111101101101000110110000000000110110000101110110101101000110110000000000110110000101101000000110110000101110110000101101000110110000101101101110110000000000110110000101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101110110000101101101101110110000101110110000101101101110110000101101101110110000101101110110110101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101101110110110110000101110110000101110110000101101101110110000101101101110110000101101110110110110110110000101101111000000111101101101101110110000101101110110110110110110000101101110110000101101101101000000110110000110110000101110110000101101101110110000101101101110110000101101110110000110110110000101101111000000111101101101101110110000101101110110000000110110000101101110110000101101101101101101110110000110110000101110110000101101101110110000101101101110110000101101110110000000110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101110110101101110110000110110110110110110000110110101110110000101110110110110110110000110110000101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101101110110110110000000101110110110110000000101110110110000000101110110110110110110000110110000101101110000101101111000000111101101101101101000000101101101000000101101000000101101101000000101101101101000000000000101101101000000000000101101101000000000101101101000000000000000000101000000101101101000101101111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam start_scene_map_on  = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111101101110110110110110110101101101110110101101101110110110110110110101101110110110110101101110110101101110110101101110110110110110101110110110110110110101110101101101110110101101101111000000111101101110110110110110110000101110000000110101101110110110110110110000110110000000110110101110110000101110110000101110110110110000000110110110110110110000110110101101110110000101101111000000111101101101000110110000000000110110000101110110101101000110110000000000110110000101101000000110110000101110110000101101000110110000101101101110110000000000110110000101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101110110000101101101101110110000101110110000101101101110110000101101101110110000101101110110110101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101101110110110110000101110110000101110110000101101101110110000101101101110110000101101110110110110110110000101101111000000111101101101101110110000101101110110110110110110000101101110110000101101101101000000110110000110110000101110110000101101101110110000101101101110110000101101110110000110110110000101101111000000111101101101101110110000101101110110000000110110000101101110110000101101101101101101110110000110110000101110110000101101101110110000101101101110110000101101110110000000110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101110110101101110110000110110110110110110000110110101110110000101110110110110110110000110110000101110110000101101111000000111101101101101110110000101101110110000101110110000101101110110000101101101110110110110000000101110110110110000000101110110110000000101110110110110110110000110110000101101110000101101111000000111101101101101101000000101101101000000101101000000101101101000000101101101101000000000000101101101000000000000101101101000000000101101101000000000000000000101000000101101101000101101111000000111101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101101111000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000000000111000000111000000111000111000111000000000111111000000111000111000111111111000111111111000111111111000111000000111000000000111000111000111000111000111000000000111000000000111000000000000000111000111000111111000111000111000111000000000111000111000111000111000000111000000000111000000111000111000111111000111000000000111111111000111111111000111111111000111111111000111111111000000000111111111000111000111111000000111000000000000111111000000111000111000000111000000000111000000111000111000111000111111000000000111000000000111111000000111000000000000000111000000000111000000000111000111000111000000111000000111000000000000111000111000111000111000000111000000000111000000111000111000111000000111000000000111000000000111000111000111111111000111111111000111111111000000000111000111000111000000111000000111000000000000111111000000111111111000000111000000000111000000111111111000111000000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam empty_on            = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000111111111111000000000000000000000111111111111000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000000000000000000000000000000111111111111000000000000000000000111111111111000000000000000000000000000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000000000000000000000000000111111111111111000000000000000000111111111111000000000000000000000000000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000000000000000000000000000111111111111111000000000000000000111111111111000000000000000000000000000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000111111111111000000000000000111111111111111000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam empty_off           = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam rickroll_on         = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111111111000111111111000111111111000111000111000000000000111111111000111111111000111000000000111000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000111000111000000111000000111000000000111000111000000000000111000111000111000111000111000000000111000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000111111111000000111000000111000000000111111000000000000000111111111000111000111000111000000000111000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000111111000000000111000000111000000000111000111000000000000111111000000111000111000111000000000111000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000111000111000111111111000111111111000111000111000000000000111000111000111111111000111111111000111111111000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam rickroll_off        = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111111111000111111111000111111111000111000111000000000000111111111000111111111000111000000000111000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000111000111000000111000000111000000000111000111000000000000111000111000111000111000111000000000111000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000111111111000000111000000111000000000111111000000000000000111111111000111000111000111000000000111000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000111111000000000111000000111000000000111000111000000000000111111000000111000111000111000000000111000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000111000111000111111111000111111111000111000111000000000000111000111000111111111000111111111000111111111000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam yareyare_on         = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111000111000000111000000111111111000111111111000000000000111000111000000111000000111111111000111111111000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000111000111000111000111000111000111000111000000000000000000111000111000111000111000111000111000111000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000111000000111111111000111111111000111111111000000000000000111000000111111111000111111111000111111111000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000111000000111000111000111111000000111000000000000000000000111000000111000111000111111000000111000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000111000000111000111000111000111000111111111000000000000000111000000111000111000111000111000111111111000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam yareyare_off        = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000111000111000000111000000111111111000111111111000000000000111000111000000111000000111111111000111111111000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000111000111000111000111000111000111000111000000000000000000111000111000111000111000111000111000111000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000111000000111111111000111111111000111111111000000000000000111000000111111111000111111111000111111111000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000111000000111000111000111111000000111000000000000000000000111000000111000111000111111000000111000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000111000000111000111000111000111000111111111000000000000000111000000111000111000111000111000111111111000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam maddeo_on           = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000111000111000000000111000000111111000000111111000000111111111000111111111000000000000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000000000000000111000111000111000111000111000111000111000111000111000111000000000111000111000000000000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000000000000111000000000111000111111111000111000111000111000111000111111111000111000111000000000000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000000000000111000000000111000111000111000111000111000111000111000111000000000111000111000000000000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000000000000111000000000111000111000111000111111000000111111000000111111111000111111111000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111110110110111111000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    localparam maddeo_off          = 6144'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111111111000111111111000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000111000000000111000000000111000000000111000000000111000000000000111000000000000000111000000000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000000000111111111000111111111000111000000000111111111000111000000000000111000000000000000111111111000111000111000111000111000111000111000111111111000000000000000000000000000000000000000000000000000000000000111000111000000000111000000000111000000000111000000000000111000000000000000000000111000111000111000111000111000111000111000000000111000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000111000000000000000111111111000111111111000111000111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000111000111000000000111000000111111000000111111000000111111111000111111111000000000000000000000111111111111111111111111000000000000000000000000000000000000111100111111000000000000000000000000111000111000111000111000111000111000111000111000111000111000000000111000111000000000000000000000111001001001001001111111000000000000000000000000000000000111100100100111111000000000000000000000111000000000111000111111111000111000111000111000111000111111111000111000111000000000000000000000000111001001001111111000000000000000000000000000000000111100100100100100111111000000000000000000111000000000111000111000111000111000111000111000111000111000000000111000111000000000000000000000000000111001111111000000000000000000000000000000000000111111111111111111111111000000000000000000111000000000111000111000111000111111000000111111000000111111111000111111111000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111111111000111111111000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111111111000111000111000000111000000111111111000111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110110110000000000000111000000000111000111000000111000000111000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111000111000111000000111000000111111111000111000111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    // State transition logic
    always @(posedge clk or posedge rst) begin
        if (rst) begin
            menuMap <= start_scene_map_off;
            counter <= 0;
            toggle <= 0;
        end else begin
            case (current_state)
                START_SCENE: begin
                    counter <= counter + 1'd1;
                    if (counter == animation_fps) begin
                        toggle <= ~toggle;
                        counter <= 0;
                    end
                    if (toggle) begin
                        menuMap <= start_scene_map_on;
                    end else begin
                        menuMap <= start_scene_map_off;
                    end
                end
                SONG_SELECT: begin
                    case (selected_song)
                        2'd0: begin // empty select
                            counter <= counter + 1'd1;
                            if (counter == animation_fps) begin
                                toggle <= ~toggle;
                                counter <= 0;
                            end
                            if (toggle) begin
                                menuMap <= empty_on;
                            end else begin
                                menuMap <= empty_off;
                            end  
                        end
                        2'd1: begin // rick roll
                            counter <= counter + 1'd1;
                            if (counter == animation_fps) begin
                                toggle <= ~toggle;
                                counter <= 0;
                            end
                            if (toggle) begin
                                menuMap <= rickroll_on;
                            end else begin
                                menuMap <= rickroll_off;
                            end  
                        end
                        2'd2: begin // Yare Yare
                            counter <= counter + 1'd1;
                            if (counter == animation_fps) begin
                                toggle <= ~toggle;
                                counter <= 0;
                            end
                            if (toggle) begin
                                menuMap <= yareyare_on;
                            end else begin
                                menuMap <= yareyare_off;
                            end  
                        end
                        2'd3: begin // Maddeo
                            counter <= counter + 1'd1;
                            if (counter == animation_fps) begin
                                toggle <= ~toggle;
                                counter <= 0;
                            end
                            if (toggle) begin
                                menuMap <= maddeo_on;
                            end else begin
                                menuMap <= maddeo_off;
                            end  
                        end
                    endcase
                end
                GAME_PLAY: begin
                    menuMap <= 0;
                end
                GAME_OVER: begin
                    menuMap <= 0;
                end
                default: begin
                    menuMap <= rickroll_on;
                end
            endcase
        end
    end
endmodule